`include "mul2.v"

module mul2tb();

endmodule