module mul2(input a,output y);

endmodule