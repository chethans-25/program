module hello;
initial
begin
$display("Hello worldd");
end
endmodule